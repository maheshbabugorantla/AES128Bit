// $Id: $
// File name:   encryption_controller.sv
// Created:     3/15/2017
// Author:      Mahesh Babu Gorantla
// Lab Section: 337-02
// Version:     1.0  Initial Design Entry
// Description: "This the main controller to orchestrate all the operations to peform the AES 128 Bit Encryption Block"
