// $Id: $
// File name:   roundKey.sv
// Created:     3/14/2017
// Author:      Mahesh Babu Gorantla
// Lab Section: 337-02
// Version:     1.0  Initial Design Entry
// Description: "This module is used to generate an individual round key for the Key Schedule"

module roundKey
(
	input wire [127:0] inputKey,
	input wire [3:0] count,
	output wire [127:0] outputRoundKey
);

	
	

endmodule 