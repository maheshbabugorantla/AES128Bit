// $Id: $
// File name:   mix_columns.sv
// Created:     3/12/2017
// Author:      Mahesh Babu Gorantla
// Lab Section: 337-02
// Version:     1.0  Initial Design Entry
// Description: "This module is used to perform the mix columns section of the AES Encryption"

module mix_columns
(
	input wire [127:0] dataIn,
	output wire [127:0] dataOut
);

	

endmodule 