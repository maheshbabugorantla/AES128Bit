// $Id: $
// File name:   decryption_block.sv
// Created:     3/17/2017
// Author:      Mahesh Babu Gorantla
// Lab Section: 337-02
// Version:     1.0  Initial Design Entry
// Description: "This is a top-level module for the AES 128-Bit Decryption Block"

module decryption_block
(
	input wire
);

endmodule 