// $Id: $
// File name:   sbox_unit.sv
// Created:     2/8/2017
// Author:      Mahesh Babu Gorantla
// Lab Section: 337-02
// Version:     1.0  Initial Design Entry
// Description: "This acts as an individual unit to the SBox"

module sbox_unit
(
	input wire [7:0] dataIn,
	output reg [7:0] byteSOut
);
	
	always_comb
	begin
		case(dataIn)
			8'h00: begin byteSOut = 8'h63; end
			8'h01: begin byteSOut = 8'h7C; end
			8'h02: begin byteSOut = 8'h77; end
			8'h03: begin byteSOut = 8'h7B; end
			8'h04: begin byteSOut = 8'hF2; end
			8'h05: begin byteSOut = 8'h6B; end
			8'h06: begin byteSOut = 8'h6F; end
			8'h07: begin byteSOut = 8'hC5; end
			8'h08: begin byteSOut = 8'h30; end
			8'h09: begin byteSOut = 8'h01; end
			8'h0A: begin byteSOut = 8'h67; end
			8'h0B: begin byteSOut = 8'h2B; end
			8'h0C: begin byteSOut = 8'hFE; end
			8'h0D: begin byteSOut = 8'hD7; end
			8'h0E: begin byteSOut = 8'hAB; end
			8'h0F: begin byteSOut = 8'h76; end
			8'h10: begin byteSOut = 8'hCA; end
			8'h11: begin byteSOut = 8'h82; end
			8'h12: begin byteSOut = 8'hC9; end
			8'h13: begin byteSOut = 8'h7D; end
			8'h14: begin byteSOut = 8'hFA; end
			8'h15: begin byteSOut = 8'h59; end
			8'h16: begin byteSOut = 8'h47; end
			8'h17: begin byteSOut = 8'hF0; end
			8'h18: begin byteSOut = 8'hAD; end
			8'h19: begin byteSOut = 8'hD4; end
			8'h1A: begin byteSOut = 8'hA2; end
			8'h1B: begin byteSOut = 8'hAF; end
			8'h1C: begin byteSOut = 8'h9C; end
			8'h1D: begin byteSOut = 8'hA4; end
			8'h1E: begin byteSOut = 8'h72; end
			8'h1F: begin byteSOut = 8'hC0; end
			8'h20: begin byteSOut = 8'hB7; end
			8'h21: begin byteSOut = 8'hFD; end
			8'h22: begin byteSOut = 8'h93; end
			8'h23: begin byteSOut = 8'h26; end
			8'h24: begin byteSOut = 8'h36; end
			8'h25: begin byteSOut = 8'h3F; end
			8'h26: begin byteSOut = 8'hF7; end
			8'h27: begin byteSOut = 8'hCC; end
			8'h28: begin byteSOut = 8'h34; end
			8'h29: begin byteSOut = 8'hA5; end
			8'h2A: begin byteSOut = 8'hE5; end
			8'h2B: begin byteSOut = 8'hF1; end
			8'h2C: begin byteSOut = 8'h71; end
			8'h2D: begin byteSOut = 8'hD8; end
			8'h2E: begin byteSOut = 8'h31; end
			8'h2F: begin byteSOut = 8'h15; end
			8'h30: begin byteSOut = 8'h04; end
			8'h31: begin byteSOut = 8'hC7; end
			8'h32: begin byteSOut = 8'h23; end
			8'h33: begin byteSOut = 8'hC3; end
			8'h34: begin byteSOut = 8'h18; end
			8'h35: begin byteSOut = 8'h96; end
			8'h36: begin byteSOut = 8'h05; end
			8'h37: begin byteSOut = 8'h9A; end
			8'h38: begin byteSOut = 8'h07; end
			8'h39: begin byteSOut = 8'h12; end
			8'h3A: begin byteSOut = 8'h80; end
			8'h3B: begin byteSOut = 8'hE2; end
			8'h3C: begin byteSOut = 8'hEB; end
			8'h3D: begin byteSOut = 8'h27; end
			8'h3E: begin byteSOut = 8'hB2; end
			8'h3F: begin byteSOut = 8'h75; end
			8'h40: begin byteSOut = 8'h09; end
			8'h41: begin byteSOut = 8'h83; end
			8'h42: begin byteSOut = 8'h2C; end
			8'h43: begin byteSOut = 8'h1A; end
			8'h44: begin byteSOut = 8'h1B; end
			8'h45: begin byteSOut = 8'h6E; end
			8'h46: begin byteSOut = 8'h5A; end
			8'h47: begin byteSOut = 8'hA0; end
			8'h48: begin byteSOut = 8'h52; end
			8'h49: begin byteSOut = 8'h3B; end
			8'h4A: begin byteSOut = 8'hD6; end
			8'h4B: begin byteSOut = 8'hB3; end
			8'h4C: begin byteSOut = 8'h29; end
			8'h4D: begin byteSOut = 8'hE3; end
			8'h4E: begin byteSOut = 8'h2F; end
			8'h4F: begin byteSOut = 8'h84; end
			8'h50: begin byteSOut = 8'h53; end
			8'h51: begin byteSOut = 8'hD1; end
			8'h52: begin byteSOut = 8'h00; end
			8'h53: begin byteSOut = 8'hED; end
			8'h54: begin byteSOut = 8'h20; end
			8'h55: begin byteSOut = 8'hFC; end
			8'h56: begin byteSOut = 8'hB1; end
			8'h57: begin byteSOut = 8'h5B; end
			8'h58: begin byteSOut = 8'h6A; end
			8'h59: begin byteSOut = 8'hCB; end
			8'h5A: begin byteSOut = 8'hBE; end
			8'h5B: begin byteSOut = 8'h39; end
			8'h5C: begin byteSOut = 8'h4A; end
			8'h5D: begin byteSOut = 8'h4C; end
			8'h5E: begin byteSOut = 8'h58; end
			8'h5F: begin byteSOut = 8'hCF; end
			8'h60: begin byteSOut = 8'hD0; end
			8'h61: begin byteSOut = 8'hEF; end
			8'h62: begin byteSOut = 8'hAA; end
			8'h63: begin byteSOut = 8'hFB; end
			8'h64: begin byteSOut = 8'h43; end
			8'h65: begin byteSOut = 8'h4D; end
			8'h66: begin byteSOut = 8'h33; end
			8'h67: begin byteSOut = 8'h85; end
			8'h68: begin byteSOut = 8'h45; end
			8'h69: begin byteSOut = 8'hF9; end
			8'h6A: begin byteSOut = 8'h02; end
			8'h6B: begin byteSOut = 8'h7F; end
			8'h6C: begin byteSOut = 8'h50; end
			8'h6D: begin byteSOut = 8'h3C; end
			8'h6E: begin byteSOut = 8'h9F; end
			8'h6F: begin byteSOut = 8'hA8; end
			8'h70: begin byteSOut = 8'h51; end
			8'h71: begin byteSOut = 8'hA3; end
			8'h72: begin byteSOut = 8'h40; end
			8'h73: begin byteSOut = 8'h8F; end
			8'h74: begin byteSOut = 8'h92; end
			8'h75: begin byteSOut = 8'h9D; end
			8'h76: begin byteSOut = 8'h38; end
			8'h77: begin byteSOut = 8'hF5; end
			8'h78: begin byteSOut = 8'hBC; end
			8'h79: begin byteSOut = 8'hB6; end
			8'h7A: begin byteSOut = 8'hDA; end
			8'h7B: begin byteSOut = 8'h21; end
			8'h7C: begin byteSOut = 8'h10; end
			8'h7D: begin byteSOut = 8'hFF; end
			8'h7E: begin byteSOut = 8'hF3; end
			8'h7F: begin byteSOut = 8'hD2; end
			8'h80: begin byteSOut = 8'hCD; end
			8'h81: begin byteSOut = 8'h0C; end
			8'h82: begin byteSOut = 8'h13; end
			8'h83: begin byteSOut = 8'hEC; end
			8'h84: begin byteSOut = 8'h5F; end
			8'h85: begin byteSOut = 8'h97; end
			8'h86: begin byteSOut = 8'h44; end
			8'h87: begin byteSOut = 8'h17; end
			8'h88: begin byteSOut = 8'hC4; end
			8'h89: begin byteSOut = 8'hA7; end
			8'h8A: begin byteSOut = 8'h7E; end
			8'h8B: begin byteSOut = 8'h3D; end
			8'h8C: begin byteSOut = 8'h64; end
			8'h8D: begin byteSOut = 8'h5D; end
			8'h8E: begin byteSOut = 8'h19; end
			8'h8F: begin byteSOut = 8'h73; end
			8'h90: begin byteSOut = 8'h60; end
			8'h91: begin byteSOut = 8'h81; end
			8'h92: begin byteSOut = 8'h4F; end
			8'h93: begin byteSOut = 8'hDC; end
			8'h94: begin byteSOut = 8'h22; end
			8'h95: begin byteSOut = 8'h2A; end
			8'h96: begin byteSOut = 8'h90; end
			8'h97: begin byteSOut = 8'h88; end
			8'h98: begin byteSOut = 8'h46; end
			8'h99: begin byteSOut = 8'hEE; end
			8'h9A: begin byteSOut = 8'hB8; end
			8'h9B: begin byteSOut = 8'h14; end
			8'h9C: begin byteSOut = 8'hDE; end
			8'h9D: begin byteSOut = 8'h5E; end
			8'h9E: begin byteSOut = 8'h0B; end
			8'h9F: begin byteSOut = 8'hDB; end
			8'hA0: begin byteSOut = 8'hE0; end
			8'hA1: begin byteSOut = 8'h32; end
			8'hA2: begin byteSOut = 8'h3A; end
			8'hA3: begin byteSOut = 8'h0A; end
			8'hA4: begin byteSOut = 8'h49; end
			8'hA5: begin byteSOut = 8'h06; end
			8'hA6: begin byteSOut = 8'h24; end
			8'hA7: begin byteSOut = 8'h5C; end
			8'hA8: begin byteSOut = 8'hC2; end
			8'hA9: begin byteSOut = 8'hD3; end
			8'hAA: begin byteSOut = 8'hAC; end
			8'hAB: begin byteSOut = 8'h62; end
			8'hAC: begin byteSOut = 8'h91; end
			8'hAD: begin byteSOut = 8'h95; end
			8'hAE: begin byteSOut = 8'hE4; end
			8'hAF: begin byteSOut = 8'h79; end
			8'hB0: begin byteSOut = 8'hE7; end
			8'hB1: begin byteSOut = 8'hC8; end
			8'hB2: begin byteSOut = 8'h37; end
			8'hB3: begin byteSOut = 8'h6D; end
			8'hB4: begin byteSOut = 8'h8D; end
			8'hB5: begin byteSOut = 8'hD5; end
			8'hB6: begin byteSOut = 8'h4E; end
			8'hB7: begin byteSOut = 8'hA9; end
			8'hB8: begin byteSOut = 8'h6C; end
			8'hB9: begin byteSOut = 8'h56; end
			8'hBA: begin byteSOut = 8'hF4; end
			8'hBB: begin byteSOut = 8'hEA; end
			8'hBC: begin byteSOut = 8'h65; end
			8'hBD: begin byteSOut = 8'h7A; end
			8'hBE: begin byteSOut = 8'hAE; end
			8'hBF: begin byteSOut = 8'h08; end
			8'hC0: begin byteSOut = 8'hBA; end
			8'hC1: begin byteSOut = 8'h78; end
			8'hC2: begin byteSOut = 8'h25; end
			8'hC3: begin byteSOut = 8'h2E; end
			8'hC4: begin byteSOut = 8'h1C; end
			8'hC5: begin byteSOut = 8'hA6; end
			8'hC6: begin byteSOut = 8'hB4; end
			8'hC7: begin byteSOut = 8'hC6; end
			8'hC8: begin byteSOut = 8'hE8; end
			8'hC9: begin byteSOut = 8'hDD; end
			8'hCA: begin byteSOut = 8'h74; end
			8'hCB: begin byteSOut = 8'h1F; end
			8'hCC: begin byteSOut = 8'h4B; end
			8'hCD: begin byteSOut = 8'hBD; end
			8'hCE: begin byteSOut = 8'h8B; end
			8'hCF: begin byteSOut = 8'h8A; end
			8'hD0: begin byteSOut = 8'h70; end
			8'hD1: begin byteSOut = 8'h3E; end
			8'hD2: begin byteSOut = 8'hB5; end
			8'hD3: begin byteSOut = 8'h66; end
			8'hD4: begin byteSOut = 8'h48; end
			8'hD5: begin byteSOut = 8'h03; end
			8'hD6: begin byteSOut = 8'hF6; end
			8'hD7: begin byteSOut = 8'h0E; end
			8'hD8: begin byteSOut = 8'h61; end
			8'hD9: begin byteSOut = 8'h35; end
			8'hDA: begin byteSOut = 8'h57; end
			8'hDB: begin byteSOut = 8'hB9; end
			8'hDC: begin byteSOut = 8'h86; end
			8'hDD: begin byteSOut = 8'hC1; end
			8'hDE: begin byteSOut = 8'h1D; end
			8'hDF: begin byteSOut = 8'h9E; end
			8'hE0: begin byteSOut = 8'hE1; end
			8'hE1: begin byteSOut = 8'hF8; end
			8'hE2: begin byteSOut = 8'h98; end
			8'hE3: begin byteSOut = 8'h11; end
			8'hE4: begin byteSOut = 8'h69; end
			8'hE5: begin byteSOut = 8'hD9; end
			8'hE6: begin byteSOut = 8'h8E; end
			8'hE7: begin byteSOut = 8'h94; end
			8'hE8: begin byteSOut = 8'h9B; end
			8'hE9: begin byteSOut = 8'h1E; end
			8'hEA: begin byteSOut = 8'h87; end
			8'hEB: begin byteSOut = 8'hE9; end
			8'hEC: begin byteSOut = 8'hCE; end
			8'hED: begin byteSOut = 8'h55; end
			8'hEE: begin byteSOut = 8'h28; end
			8'hEF: begin byteSOut = 8'hDF; end
			8'hF0: begin byteSOut = 8'h8C; end
			8'hF1: begin byteSOut = 8'hA1; end
			8'hF2: begin byteSOut = 8'h89; end
			8'hF3: begin byteSOut = 8'h0D; end
			8'hF4: begin byteSOut = 8'hBF; end
			8'hF5: begin byteSOut = 8'hE6; end
			8'hF6: begin byteSOut = 8'h42; end
			8'hF7: begin byteSOut = 8'h68; end
			8'hF8: begin byteSOut = 8'h41; end
			8'hF9: begin byteSOut = 8'h99; end
			8'hFA: begin byteSOut = 8'h2D; end
			8'hFB: begin byteSOut = 8'h0F; end
			8'hFC: begin byteSOut = 8'hB0; end
			8'hFD: begin byteSOut = 8'h54; end
			8'hFE: begin byteSOut = 8'hBB; end
			8'hFF: begin byteSOut = 8'h16; end
			default: begin byteSOut = 8'h00; end
		endcase
	end

endmodule 