// $Id: $
// File name:   tb_KeySchedule.sv
// Created:     3/14/2017
// Author:      Mahesh Babu Gorantla
// Lab Section: 337-02
// Version:     1.0  Initial Design Entry
// Description: This is the testbench to test the proper working of the KeySchedule for the 128-bit Key Schedule
