// $Id: $
// File name:   top_level_controller.sv
// Created:     4/11/2017
// Author:      Mahesh Babu Gorantla
// Lab Section: 337-02
// Version:     1.0  Initial Design Entry
// Description: "This is the Main Controller for the Top-Level Block for the Project"
