// $Id: $
// File name:   tb_decryption_controller.sv
// Created:     3/15/2017
// Author:      Mahesh Babu Gorantla
// Lab Section: 337-02
// Version:     1.0  Initial Design Entry
// Description: 
// "This is the testbench for decryption_controller"
