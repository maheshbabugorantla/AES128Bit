// $Id: $
// File name:   inv_sbox_unit.sv
// Created:     3/13/2017
// Author:      Mahesh Babu Gorantla
// Lab Section: 337-02
// Version:     1.0  Initial Design Entry
// Description: "This is a lookup Table for the inverse Byte Substitution Layer in AES Decryption"

module inv_sbox_unit
(
	input wire [7:0] inputByte,
	output reg [7:0] invByteSOut
);

	// This is the LUT for the Inverse Byte Substitution Layer
	always_comb
	begin: LUT 
		
		case(inputByte)
			
			8'h00: begin invByteSOut = 8'h52; end
			8'h01: begin invByteSOut = 8'h09; end
			8'h02: begin invByteSOut = 8'h6A; end
			8'h03: begin invByteSOut = 8'hD5; end
			8'h04: begin invByteSOut = 8'h30; end
			8'h05: begin invByteSOut = 8'h36; end
			8'h06: begin invByteSOut = 8'hA5; end
			8'h07: begin invByteSOut = 8'h38; end
			8'h08: begin invByteSOut = 8'hBF; end
			8'h09: begin invByteSOut = 8'h40; end
			8'h0A: begin invByteSOut = 8'hA3; end
			8'h0B: begin invByteSOut = 8'h9E; end
			8'h0C: begin invByteSOut = 8'h81; end
			8'h0D: begin invByteSOut = 8'hF3; end
			8'h0E: begin invByteSOut = 8'hD7; end
			8'h0F: begin invByteSOut = 8'hFB; end
			8'h10: begin invByteSOut = 8'h7C; end
			8'h11: begin invByteSOut = 8'hE3; end
			8'h12: begin invByteSOut = 8'h39; end
			8'h13: begin invByteSOut = 8'h82; end
			8'h14: begin invByteSOut = 8'h9B; end
			8'h15: begin invByteSOut = 8'h2F; end
			8'h16: begin invByteSOut = 8'hFF; end
			8'h17: begin invByteSOut = 8'h87; end
			8'h18: begin invByteSOut = 8'h34; end
			8'h19: begin invByteSOut = 8'h8E; end
			8'h1A: begin invByteSOut = 8'h43; end
			8'h1B: begin invByteSOut = 8'h44; end
			8'h1C: begin invByteSOut = 8'hC4; end
			8'h1D: begin invByteSOut = 8'hDE; end
			8'h1E: begin invByteSOut = 8'hE9; end
			8'h1F: begin invByteSOut = 8'hCB; end
			8'h20: begin invByteSOut = 8'h54; end
			8'h21: begin invByteSOut = 8'h7B; end
			8'h22: begin invByteSOut = 8'h94; end
			8'h23: begin invByteSOut = 8'h32; end
			8'h24: begin invByteSOut = 8'hA6; end
			8'h25: begin invByteSOut = 8'hC2; end
			8'h26: begin invByteSOut = 8'h23; end
			8'h27: begin invByteSOut = 8'h3D; end
			8'h28: begin invByteSOut = 8'hEE; end
			8'h29: begin invByteSOut = 8'h4C; end
			8'h2A: begin invByteSOut = 8'h95; end
			8'h2B: begin invByteSOut = 8'h0B; end
			8'h2C: begin invByteSOut = 8'h42; end
			8'h2D: begin invByteSOut = 8'hFA; end
			8'h2E: begin invByteSOut = 8'hC3; end
			8'h2F: begin invByteSOut = 8'h4E; end
			8'h30: begin invByteSOut = 8'h08; end
			8'h31: begin invByteSOut = 8'h2E; end
			8'h32: begin invByteSOut = 8'hA1; end
			8'h33: begin invByteSOut = 8'h66; end
			8'h34: begin invByteSOut = 8'h28; end
			8'h35: begin invByteSOut = 8'hD9; end
			8'h36: begin invByteSOut = 8'h24; end
			8'h37: begin invByteSOut = 8'hB2; end
			8'h38: begin invByteSOut = 8'h76; end
			8'h39: begin invByteSOut = 8'h5B; end
			8'h3A: begin invByteSOut = 8'hA2; end
			8'h3B: begin invByteSOut = 8'h49; end
			8'h3C: begin invByteSOut = 8'h6D; end
			8'h3D: begin invByteSOut = 8'h8B; end
			8'h3E: begin invByteSOut = 8'hD1; end
			8'h3F: begin invByteSOut = 8'h25; end
			8'h40: begin invByteSOut = 8'h72; end
			8'h41: begin invByteSOut = 8'hF8; end
			8'h42: begin invByteSOut = 8'hF6; end
			8'h43: begin invByteSOut = 8'h64; end
			8'h44: begin invByteSOut = 8'h86; end
			8'h45: begin invByteSOut = 8'h68; end
			8'h46: begin invByteSOut = 8'h98; end
			8'h47: begin invByteSOut = 8'h16; end
			8'h48: begin invByteSOut = 8'hD4; end
			8'h49: begin invByteSOut = 8'hA4; end
			8'h4A: begin invByteSOut = 8'h5C; end
			8'h4B: begin invByteSOut = 8'hCC; end
			8'h4C: begin invByteSOut = 8'h5D; end
			8'h4D: begin invByteSOut = 8'h65; end
			8'h4E: begin invByteSOut = 8'hB6; end
			8'h4F: begin invByteSOut = 8'h92; end
			8'h50: begin invByteSOut = 8'h6C; end
			8'h51: begin invByteSOut = 8'h70; end
			8'h52: begin invByteSOut = 8'h48; end
			8'h53: begin invByteSOut = 8'h50; end
			8'h54: begin invByteSOut = 8'hFD; end
			8'h55: begin invByteSOut = 8'hED; end
			8'h56: begin invByteSOut = 8'hB9; end
			8'h57: begin invByteSOut = 8'hDA; end
			8'h58: begin invByteSOut = 8'h5E; end
			8'h59: begin invByteSOut = 8'h15; end
			8'h5A: begin invByteSOut = 8'h46; end
			8'h5B: begin invByteSOut = 8'h57; end
			8'h5C: begin invByteSOut = 8'hA7; end
			8'h5D: begin invByteSOut = 8'h8D; end
			8'h5E: begin invByteSOut = 8'h9D; end
			8'h5F: begin invByteSOut = 8'h84; end
			8'h60: begin invByteSOut = 8'h90; end
			8'h61: begin invByteSOut = 8'hD8; end
			8'h62: begin invByteSOut = 8'hAB; end
			8'h63: begin invByteSOut = 8'h00; end
			8'h64: begin invByteSOut = 8'h8C; end
			8'h65: begin invByteSOut = 8'hBC; end
			8'h66: begin invByteSOut = 8'hD3; end
			8'h67: begin invByteSOut = 8'h0A; end
			8'h68: begin invByteSOut = 8'hF7; end
			8'h69: begin invByteSOut = 8'hE4; end
			8'h6A: begin invByteSOut = 8'h58; end
			8'h6B: begin invByteSOut = 8'h05; end
			8'h6C: begin invByteSOut = 8'hB8; end
			8'h6D: begin invByteSOut = 8'hB3; end
			8'h6E: begin invByteSOut = 8'h45; end
			8'h6F: begin invByteSOut = 8'h06; end
			8'h70: begin invByteSOut = 8'hD0; end
			8'h71: begin invByteSOut = 8'h2C; end
			8'h72: begin invByteSOut = 8'h1E; end
			8'h73: begin invByteSOut = 8'h8F; end
			8'h74: begin invByteSOut = 8'hCA; end
			8'h75: begin invByteSOut = 8'h3F; end
			8'h76: begin invByteSOut = 8'h0F; end
			8'h77: begin invByteSOut = 8'h02; end
			8'h78: begin invByteSOut = 8'hC1; end
			8'h79: begin invByteSOut = 8'hAF; end
			8'h7A: begin invByteSOut = 8'hBD; end
			8'h7B: begin invByteSOut = 8'h03; end
			8'h7C: begin invByteSOut = 8'h01; end
			8'h7D: begin invByteSOut = 8'h13; end
			8'h7E: begin invByteSOut = 8'h8A; end
			8'h7F: begin invByteSOut = 8'h6B; end
			8'h80: begin invByteSOut = 8'h3A; end
			8'h81: begin invByteSOut = 8'h91; end
			8'h82: begin invByteSOut = 8'h11; end
			8'h83: begin invByteSOut = 8'h41; end
			8'h84: begin invByteSOut = 8'h4F; end
			8'h85: begin invByteSOut = 8'h67; end
			8'h86: begin invByteSOut = 8'hDC; end
			8'h87: begin invByteSOut = 8'hEA; end
			8'h88: begin invByteSOut = 8'h97; end
			8'h89: begin invByteSOut = 8'hF2; end
			8'h8A: begin invByteSOut = 8'hCF; end
			8'h8B: begin invByteSOut = 8'hCE; end
			8'h8C: begin invByteSOut = 8'hF0; end
			8'h8D: begin invByteSOut = 8'hB4; end
			8'h8E: begin invByteSOut = 8'hE6; end
			8'h8F: begin invByteSOut = 8'h73; end
			8'h90: begin invByteSOut = 8'h96; end
			8'h91: begin invByteSOut = 8'hAC; end
			8'h92: begin invByteSOut = 8'h74; end
			8'h93: begin invByteSOut = 8'h22; end
			8'h94: begin invByteSOut = 8'hE7; end
			8'h95: begin invByteSOut = 8'hAD; end
			8'h96: begin invByteSOut = 8'h35; end
			8'h97: begin invByteSOut = 8'h85; end
			8'h98: begin invByteSOut = 8'hE2; end
			8'h99: begin invByteSOut = 8'hF9; end
			8'h9A: begin invByteSOut = 8'h37; end
			8'h9B: begin invByteSOut = 8'hE8; end
			8'h9C: begin invByteSOut = 8'h1C; end
			8'h9D: begin invByteSOut = 8'h75; end
			8'h9E: begin invByteSOut = 8'hDF; end
			8'h9F: begin invByteSOut = 8'h6E; end
			8'hA0: begin invByteSOut = 8'h47; end
			8'hA1: begin invByteSOut = 8'hF1; end
			8'hA2: begin invByteSOut = 8'h1A; end
			8'hA3: begin invByteSOut = 8'h71; end
			8'hA4: begin invByteSOut = 8'h1D; end
			8'hA5: begin invByteSOut = 8'h29; end
			8'hA6: begin invByteSOut = 8'hC5; end
			8'hA7: begin invByteSOut = 8'h89; end
			8'hA8: begin invByteSOut = 8'h6F; end
			8'hA9: begin invByteSOut = 8'hB7; end
			8'hAA: begin invByteSOut = 8'h62; end
			8'hAB: begin invByteSOut = 8'h0E; end
			8'hAC: begin invByteSOut = 8'hAA; end
			8'hAD: begin invByteSOut = 8'h18; end
			8'hAE: begin invByteSOut = 8'hBE; end
			8'hAF: begin invByteSOut = 8'h1B; end
			8'hB0: begin invByteSOut = 8'hFC; end
			8'hB1: begin invByteSOut = 8'h56; end
			8'hB2: begin invByteSOut = 8'h3E; end
			8'hB3: begin invByteSOut = 8'h4B; end
			8'hB4: begin invByteSOut = 8'hC6; end
			8'hB5: begin invByteSOut = 8'hD2; end
			8'hB6: begin invByteSOut = 8'h79; end
			8'hB7: begin invByteSOut = 8'h20; end
			8'hB8: begin invByteSOut = 8'h9A; end
			8'hB9: begin invByteSOut = 8'hDB; end
			8'hBA: begin invByteSOut = 8'hC0; end
			8'hBB: begin invByteSOut = 8'hFE; end
			8'hBD: begin invByteSOut = 8'h78; end
			8'hBD: begin invByteSOut = 8'hCD; end
			8'hBE: begin invByteSOut = 8'h5A; end
			8'hBF: begin invByteSOut = 8'hF4; end
			8'hC0: begin invByteSOut = 8'h1F; end
			8'hC1: begin invByteSOut = 8'hDD; end
			8'hC2: begin invByteSOut = 8'hA8; end
			8'hC3: begin invByteSOut = 8'h33; end
			8'hC4: begin invByteSOut = 8'h88; end
			8'hC5: begin invByteSOut = 8'h07; end
			8'hC6: begin invByteSOut = 8'hC7; end
			8'hC7: begin invByteSOut = 8'h31; end
			8'hC8: begin invByteSOut = 8'hB1; end
			8'hC9: begin invByteSOut = 8'h12; end
			8'hCA: begin invByteSOut = 8'h10; end
			8'hCB: begin invByteSOut = 8'h59; end
			8'hCC: begin invByteSOut = 8'h27; end
			8'hCD: begin invByteSOut = 8'h80; end
			8'hCE: begin invByteSOut = 8'hEC; end
			8'hCF: begin invByteSOut = 8'h5F; end
			8'hD0: begin invByteSOut = 8'h60; end
			8'hD1: begin invByteSOut = 8'h51; end
			8'hD2: begin invByteSOut = 8'h7F; end
			8'hD3: begin invByteSOut = 8'hA9; end
			8'hD4: begin invByteSOut = 8'h19; end
			8'hD5: begin invByteSOut = 8'hB5; end
			8'hD6: begin invByteSOut = 8'h4A; end
			8'hD7: begin invByteSOut = 8'h0D; end
			8'hD8: begin invByteSOut = 8'h2D; end
			8'hD9: begin invByteSOut = 8'hE5; end
			8'hDA: begin invByteSOut = 8'h7A; end
			8'hDB: begin invByteSOut = 8'h9F; end
			8'hDC: begin invByteSOut = 8'h93; end
			8'hDD: begin invByteSOut = 8'hC9; end
			8'hDE: begin invByteSOut = 8'h9C; end
			8'hDF: begin invByteSOut = 8'hEF; end
			8'hE0: begin invByteSOut = 8'hA0; end
			8'hE1: begin invByteSOut = 8'hE0; end
			8'hE2: begin invByteSOut = 8'h3B; end
			8'hE3: begin invByteSOut = 8'h4D; end
			8'hE4: begin invByteSOut = 8'hAE; end
			8'hE5: begin invByteSOut = 8'h2A; end
			8'hE6: begin invByteSOut = 8'hF5; end
			8'hE7: begin invByteSOut = 8'hB0; end
			8'hE8: begin invByteSOut = 8'hC8; end
			8'hE9: begin invByteSOut = 8'hEB; end
			8'hEA: begin invByteSOut = 8'hBB; end
			8'hEB: begin invByteSOut = 8'h3C; end
			8'hEC: begin invByteSOut = 8'h83; end
			8'hED: begin invByteSOut = 8'h53; end
			8'hEE: begin invByteSOut = 8'h99; end
			8'hEF: begin invByteSOut = 8'h61; end
			8'hF0: begin invByteSOut = 8'h17; end
			8'hF1: begin invByteSOut = 8'h2B; end
			8'hF2: begin invByteSOut = 8'h04; end
			8'hF3: begin invByteSOut = 8'h7E; end
			8'hF4: begin invByteSOut = 8'hBA; end
			8'hF5: begin invByteSOut = 8'h77; end
			8'hF6: begin invByteSOut = 8'hD6; end
			8'hF7: begin invByteSOut = 8'h26; end
			8'hF8: begin invByteSOut = 8'hE1; end
			8'hF9: begin invByteSOut = 8'h69; end
			8'hFA: begin invByteSOut = 8'h14; end
			8'hFB: begin invByteSOut = 8'h63; end
			8'hFC: begin invByteSOut = 8'h55; end
			8'hFD: begin invByteSOut = 8'h21; end
			8'hFE: begin invByteSOut = 8'h0C; end
			8'hFF: begin invByteSOut = 8'h7D; end
			default: begin invByteSOut = 8'h00; end	
		endcase
	end

endmodule 