// $Id: $
// File name:   decryption_controller.sv
// Created:     3/15/2017
// Author:      Mahesh Babu Gorantla
// Lab Section: 337-02
// Version:     1.0  Initial Design Entry
// Description: "This is the main controller to orchestrate all the operations to perform the AES 128 Bit Decryption"
