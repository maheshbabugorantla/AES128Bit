// $Id: $
// File name:   tb_inv_subBytes.sv
// Created:     3/13/2017
// Author:      Mahesh Babu Gorantla
// Lab Section: 337-02
// Version:     1.0  Initial Design Entry
// Description: "This is the testbench for the inv_subBytes.sv module"
